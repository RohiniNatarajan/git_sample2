nside index file
