inside index1.sv file

